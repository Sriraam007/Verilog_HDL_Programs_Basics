module COMP_2BIT(A,B,OUT3,OUT2,OUT1);
    input [1:0]A,B;
    output OUT3,OUT2,OUT1;
    